// Created by prof. Mingu Kang @VVIP Lab in UCSD ECE department
// Please do not spread this code without permission 
module mac (out, a, b, c);

parameter a_bw = 2;
parameter b_bw = 4;
parameter psum_bw = 16;

output signed [psum_bw-1:0] out;
input signed  [a_bw-1:0] a;  // activation
input signed  [b_bw-1:0] b;  // weight
input signed  [psum_bw-1:0] c;


wire signed [2*b_bw:0] product;
wire signed [psum_bw-1:0] psum;
wire signed [a_bw:0]   a_pad;

assign a_pad = {2'b00, a}; // force to be unsigned number
assign product = a_pad * b;

assign psum = product + c;
assign out = psum;

endmodule
