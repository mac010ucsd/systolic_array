module core;


parameter bw = 2;
parameter b_bw = 4;
parameter psum_bw = 32;
parameter col = 2;
parameter row = 2;




endmodule